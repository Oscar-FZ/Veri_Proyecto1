class scoreboard #(parameter bits = 1, parameter drvrs = 4, parameter pckg_sz = 16, parameter broadcast = {8{1'b1}});
    //Plan de ataque:
    //Agarrar el mensaje del checker
    //Calcular el retardo 
    //Meterlo a un archivo csv (Tiempo de envio, terminal de origen, terminal de destino, tiempo de recibido, retraso en el envio)

    //Definicion de variables
    bit inicio;
    string tipo_test;
    string nombre_archivo;
    int test_aleatorio;
    int cont;

    sb_pckg #(.drvrs(drvrs), .pckg_sz(pckg_sz)) transaccion_chkr;
  
    //Definicion de mailboxes
    test_type test_sb_mbx;
    sb_pckg_mbx #(.drvrs(drvrs), .pckg_sz(pckg_sz)) chkr_sb_mbx;

    function new();
        chkr_sb_mbx = new();
        test_sb_mbx = new();
        transaccion_chkr = new();
        inicio = 1;
        cont = 1;
        nombre_archivo = "Aleatorio.csv";
        tipo_test = "Aleatorio";
    endfunction

    task run();
        forever begin
            //wait(fin_test.triggered);
            if (inicio) begin
                test_sb_mbx.get(tipo_test);
                test_aleatorio = $fopen(nombre_archivo, "w");
                $fwrite(test_aleatorio, "Test: ", tipo_test, "\n");
                $fwrite(test_aleatorio, "Parametros del Ambiente\n");
                $fwrite(test_aleatorio, "Bits = %0d\n", bits);
                $fwrite(test_aleatorio, "Drivers = %0d\n", drvrs);
                $fwrite(test_aleatorio, "Tamaño del Paquete = %0d\n", pckg_sz);
                $fwrite(test_aleatorio, "Identificador de Broadcast = %b\n", broadcast);
                $fwrite(test_aleatorio, "Numero; Paquete; Estado; Dispositivo de Origen; Dispositivo Destino; Tiempo de Envio; Tiempo de Recibido; Latencia;\n");
                $fclose(test_aleatorio);
                inicio = 0;
            end

            else begin
                $display("[AQUI]");
                chkr_sb_mbx.get(transaccion_chkr);
                test_aleatorio = $fopen(nombre_archivo, "a");
                $fwrite(test_aleatorio, "%d; 0x%h; %b; %d; %d; %d; %d; %d; \n", cont, transaccion_chkr.dato_enviado, transaccion_chkr.completado, transaccion_chkr.disp_origen, transaccion_chkr.disp_destino, transaccion_chkr.tiempo_push, transaccion_chkr.tiempo_pop, transaccion_chkr.latencia);
                $fclose(test_aleatorio);
                cont += 1;
            end

            if ((chkr_sb_mbx.num() == 0) && (fin_test.triggered)) begin
                $finish;
            end
            //$display("Aqui va el resto ajaj equis de");
            //$finish;
      
        end
    endtask
endclass
